LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL; 
USE WORK.RV_PKG.ALL;

ENTITY ULA_RV IS 
	GENERIC (WSIZE : natural := 32);
	PORT (
		OPCODE : IN ULA_OP;
		A, B : IN STD_LOGIC_VECTOR(WSIZE-1 DOWNTO 0);
		Z : OUT STD_LOGIC_VECTOR(WSIZE-1 DOWNTO 0);
		ZERO : OUT STD_LOGIC);
END ULA_RV;

ARCHITECTURE ULA_ARCH OF ULA_RV IS
	
SIGNAL A32 : STD_LOGIC_VECTOR(WSIZE-1 DOWNTO 0);
BEGIN
	Z <= A32;
		
	PROCESS(A, B, OPCODE, A32)
	BEGIN
		IF (UNSIGNED(A32) = 0)
			THEN ZERO <= '1';
			ELSE ZERO <= '0';
		END IF;
		
		CASE OPCODE IS
			WHEN ADD_OP => A32 <= STD_LOGIC_VECTOR(SIGNED(A) + SIGNED(B));
			WHEN SUB_OP => A32 <= STD_LOGIC_VECTOR(SIGNED(A) - SIGNED(B));
			WHEN AND_OP => A32 <= A AND B;
			WHEN OR_OP => A32 <= A OR B;
			WHEN NOR_OP => A32 <= A NOR B;
			WHEN XOR_OP => A32 <= A XOR B;
			WHEN SLL_OP => A32 <= STD_LOGIC_VECTOR(SHIFT_LEFT(UNSIGNED(A), TO_INTEGER(UNSIGNED(B))));
			WHEN SRL_OP => A32 <= STD_LOGIC_VECTOR(SHIFT_RIGHT(UNSIGNED(A), TO_INTEGER(UNSIGNED(B))));
			WHEN SRA_OP => A32 <= STD_LOGIC_VECTOR(SHIFT_RIGHT(SIGNED(A), TO_INTEGER(UNSIGNED(B))));
			WHEN SLT_OP => IF(SIGNED(A) < SIGNED(B)) 
								THEN A32 <= X"00000001"; 
								ELSE A32 <= X"00000000"; 
								END IF;
			WHEN SLTU_OP => 	IF(UNSIGNED(A) < UNSIGNED(B)) 
									THEN A32 <= X"00000001"; 
									ELSE A32 <= X"00000000"; 
									END IF;
			WHEN SGE_OP => 	IF(SIGNED(A) >= SIGNED(B)) 
									THEN A32 <= X"00000001"; 
									ELSE A32 <= X"00000000"; 
									END IF;
			WHEN SGEU_OP => 	IF(UNSIGNED(A) >= UNSIGNED(B)) 
									THEN A32 <= X"00000001";  
									ELSE A32 <= X"00000000"; 
									END IF;
			WHEN SEQ_OP =>		IF(SIGNED(A) = SIGNED(B)) 
									THEN A32 <= X"00000001";  
									ELSE A32 <= X"00000000"; 
									END IF;
			WHEN SNE_OP => 	IF(SIGNED(A) /= SIGNED(B)) 
									THEN A32 <= X"00000001";  
									ELSE A32 <= X"00000000"; 
									END IF;
		END CASE;
	END PROCESS;
END ULA_ARCH;
